module xor_64 (x, y, z);

input [63:0] x, y;
output [63:0] z;

integer i;
for (i = 0; i < 64; i)
endmodule